library ieee;
use ieee.std_logic_1164.all;

package Common is
    type CellType is array (0 to 8, 0 to 1) of std_logic;
end package Common;

package body Common is
    
end package body Common;
